module mem_sim;
endmodule