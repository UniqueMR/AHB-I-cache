module cache_state_handler(
    input clk,
    input rst,

    output reg [1:0] state
);

always @(posedge clk or negedge rst)    begin
    
end


endmodule